module instruction_memory(address,data);

input [5:0] address;
output [31:0] data;

wire [31:0] rom [63:0];

assign rom[0] = 32'd0;
assign rom[1] = 32'd1;
assign rom[2] = 32'd2;
assign rom[3] = 32'd3;
assign rom[4] = 32'd4;
assign rom[5] = 32'd5;
assign rom[6] = 32'd6;
assign rom[7] = 32'd7;
assign rom[8] = 32'd8;
assign rom[9] = 32'd9;
assign rom[10] = 32'd10;
assign rom[11] = 32'd11;
assign rom[12] = 32'd12;
assign rom[13] = 32'd13;
assign rom[14] = 32'd14;
assign rom[15] = 32'd15;
assign rom[16] = 32'd16;
assign rom[17] = 32'd17;
assign rom[18] = 32'd18;
assign rom[19] = 32'd19;
assign rom[20] = 32'd20;
assign rom[21] = 32'd21;
assign rom[22] = 32'd22;
assign rom[23] = 32'd23;
assign rom[24] = 32'd24;
assign rom[25] = 32'd25;
assign rom[26] = 32'd26;
assign rom[27] = 32'd27;
assign rom[28] = 32'd28;
assign rom[29] = 32'd29;
assign rom[30] = 32'd30;
assign rom[31] = 32'd31;
assign rom[32] = 32'd32;
assign rom[33] = 32'd33;
assign rom[34] = 32'd34;
assign rom[35] = 32'd35;
assign rom[36] = 32'd36;
assign rom[37] = 32'd37;
assign rom[38] = 32'd38;
assign rom[39] = 32'd39;
assign rom[40] = 32'd40;
assign rom[41] = 32'd41;
assign rom[42] = 32'd42;
assign rom[43] = 32'd43;
assign rom[44] = 32'd44;
assign rom[45] = 32'd45;
assign rom[46] = 32'd46;
assign rom[47] = 32'd47;
assign rom[48] = 32'd48;
assign rom[49] = 32'd49;
assign rom[50] = 32'd50;
assign rom[51] = 32'd51;
assign rom[52] = 32'd52;
assign rom[53] = 32'd53;
assign rom[54] = 32'd54;
assign rom[55] = 32'd55;
assign rom[56] = 32'd56;
assign rom[57] = 32'd57;
assign rom[58] = 32'd58;
assign rom[59] = 32'd59;
assign rom[60] = 32'd60;
assign rom[61] = 32'd61;
assign rom[62] = 32'd62;
assign rom[63] = 32'd63;
assign data = rom[address];

endmodule
