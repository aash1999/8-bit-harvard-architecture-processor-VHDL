module instruction(Instruction_out, PCAdress);
	output reg [31:0] Instruction_out;
	input  [5:0] PCAdress;
	
	always @(*)
	begin
		case (PCAdress)
			32'd0:  Instruction_out = 32'b00000000000000000000000000001010;
			32'd1:  Instruction_out = 32'b00000000001000000000000000001111; 
			32'd2:  Instruction_out = 32'b00000000010000000000000000000011; 
			32'd3:  Instruction_out = 32'b00000000011000000000000000011001; 
			32'd4:  Instruction_out = 32'b00000000100000000000000000100000; 
			32'd5:  Instruction_out = 32'b00000000101000000000000000001100; 
			32'd6:  Instruction_out = 32'b00010011111100000000000000000001;
			32'd7:  Instruction_out = 32'b00010111111100010000000001100010;
			32'd8:  Instruction_out = 32'b00010111111100100000000010000101;
			32'd9:  Instruction_out = 32'b00010011111100110000001000010001;
			32'd10:  Instruction_out = 32'b00010011111101000000001001110010;
			//32'd11:  Instruction_out = 32'b00110000000100000000000001000001;
			//32'd12:  Instruction_out = 32'b00111010000000000000000000000001;
			//32'd13:  Instruction_out = 32'b00000011011000000000000000000010;
			//32'd14:  Instruction_out = 32'b00111110000110000000000000111011;
			//32'd15:  Instruction_out = 32'b00000100001000000000000000000010;
			//32'd16:  Instruction_out = 32'b00010000000100000000000000100010;
			//32'd17:  Instruction_out = 32'b00001100000000000000000000000001;
			//32'd18:  Instruction_out = 32'b00001000010000000000000000000000;
			//32'd19:  Instruction_out = 32'b00010010000110000000000000100010;
			//32'd18:  Instruction_out = 32'b;
			default: Instruction_out = 32'b00000000000000000000000000000000;

		endcase
	end
	endmodule 